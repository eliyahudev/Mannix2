 

//===============================================
//         Start Header Num 1
//===============================================

module MODULE_NAME_TEMPLATE
  (
   // System
   rf_clk,                        // [I] 1b gated clock 
   hw_reset_n,                 // [I] 1b Sync reset
   scan_mode,                  // [I] 1b scan mode for the reset ctrl block
   //===============================================
   //         End Header Num 1
   //===============================================
   
