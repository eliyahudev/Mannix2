`undef STD_DEFINED
module m_mx2( input A, input B, input S, output Z);

`ifdef STD_SIM
 `define STD_DEFINED
   assign Z = S ? B : A;

`elsif TSMC_65
   // /data/tsmc/65LP//dig_libs/ARM_FEONLY/arm/tsmc/cln65lp/sc9_base_rvt/r0p0/verilog/sc9_cln65lp_base_rvt.v
   // /data/tsmc/65LP//dig_libs/ARM_FEONLY/arm/tsmc/cln65lp/sc9_base_rvt/r0p0/doc/sc9_cln65lp_base_rvt_databook.pdf
 `define STD_DEFINED
 `define I_CLK_MX2 i_clk_mx2 (.Y(Z), .A(A), .B(B), .S0(S))

 `ifdef CTS_LVT
   MX2_X1B_A9TL `I_CLK_MX2;
 `else
   MX2_X1B_A9TR `I_CLK_MX2;
 `endif

 `undef I_CLK_MX2

`elsif TSMC16
   // /data/tsmc/16FF/dig_libs/TSMCHOME/digital/Front_End/verilog/tcbn16ffcllbwp16p90cpd_100a/tcbn16ffcllbwp16p90cpd.v
   // /data/tsmc/16FF/dig_libs/doc/DB_TCBN16FFCLLBWP16P90CPD_TT0P8V25C.pdf
 `define STD_DEFINED
 `define I_CLK_MX2 I_clk_mx2 (.Z(Z), .I0(A), .I1(B), .S(S))
 `ifdef CTS_ULVT
   CKMUX2D1BWP16P90CPDULVT `I_CLK_MX2;
 `elsif CTS_LVT
   CKMUX2D1BWP16P90CPDLVT `I_CLK_MX2;
 `else
   CKMUX2D1BWP16P90CPD `I_CLK_MX2;
 `endif

 `undef I_CLK_MX2

`endif // !`elsif TSMC16


endmodule
`ifndef STD_DEFINED
    ERROR NO STD_X TECHNOLOGY FOUND
`endif
