endmodule 
//==========================================
//         End Header Num 3
//==========================================



