VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO spram_1024x16m8b1pm2re1
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN spram_1024x16m8b1pm2re1 0 0 ;
  SIZE 89.774 BY 195.084 ;
  SYMMETRY X Y  ;
  PIN Q[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    ANTENNADIFFAREA 0.168 ;
    PORT
      LAYER M2 ;
        RECT 0.118 7.061 0.358 7.201 ;
    END
  END Q[0]
  PIN Q[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    ANTENNADIFFAREA 0.168 ;
    PORT
      LAYER M2 ;
        RECT 0.118 15.573 0.358 15.713 ;
    END
  END Q[1]
  PIN Q[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    ANTENNADIFFAREA 0.168 ;
    PORT
      LAYER M2 ;
        RECT 0.118 24.085 0.358 24.225 ;
    END
  END Q[2]
  PIN Q[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    ANTENNADIFFAREA 0.168 ;
    PORT
      LAYER M2 ;
        RECT 0.118 32.597 0.358 32.737 ;
    END
  END Q[3]
  PIN Q[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    ANTENNADIFFAREA 0.168 ;
    PORT
      LAYER M2 ;
        RECT 0.118 41.109 0.358 41.249 ;
    END
  END Q[4]
  PIN Q[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    ANTENNADIFFAREA 0.168 ;
    PORT
      LAYER M2 ;
        RECT 0.118 49.621 0.358 49.761 ;
    END
  END Q[5]
  PIN Q[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    ANTENNADIFFAREA 0.168 ;
    PORT
      LAYER M2 ;
        RECT 0.118 58.133 0.358 58.273 ;
    END
  END Q[6]
  PIN Q[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    ANTENNADIFFAREA 0.168 ;
    PORT
      LAYER M2 ;
        RECT 0.118 66.645 0.358 66.785 ;
    END
  END Q[7]
  PIN D[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    ANTENNADIFFAREA 0.056 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.06 ;
    PORT
      LAYER M2 ;
        RECT 0.118 5.705 0.358 5.805 ;
    END
  END D[0]
  PIN D[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    ANTENNADIFFAREA 0.056 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.06 ;
    PORT
      LAYER M2 ;
        RECT 0.118 14.217 0.358 14.317 ;
    END
  END D[1]
  PIN D[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    ANTENNADIFFAREA 0.056 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.06 ;
    PORT
      LAYER M2 ;
        RECT 0.118 22.729 0.358 22.829 ;
    END
  END D[2]
  PIN D[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    ANTENNADIFFAREA 0.056 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.06 ;
    PORT
      LAYER M2 ;
        RECT 0.118 31.241 0.358 31.341 ;
    END
  END D[3]
  PIN D[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    ANTENNADIFFAREA 0.056 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.06 ;
    PORT
      LAYER M2 ;
        RECT 0.118 39.753 0.358 39.853 ;
    END
  END D[4]
  PIN D[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    ANTENNADIFFAREA 0.056 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.06 ;
    PORT
      LAYER M2 ;
        RECT 0.118 48.265 0.358 48.365 ;
    END
  END D[5]
  PIN D[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    ANTENNADIFFAREA 0.056 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.06 ;
    PORT
      LAYER M2 ;
        RECT 0.118 56.777 0.358 56.877 ;
    END
  END D[6]
  PIN D[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    ANTENNADIFFAREA 0.056 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.06 ;
    PORT
      LAYER M2 ;
        RECT 0.118 65.289 0.358 65.389 ;
    END
  END D[7]
  PIN TD[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    ANTENNADIFFAREA 0.056 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.06 ;
    PORT
      LAYER M2 ;
        RECT 0.118 6.135 0.358 6.235 ;
    END
  END TD[0]
  PIN TD[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    ANTENNADIFFAREA 0.056 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.06 ;
    PORT
      LAYER M2 ;
        RECT 0.118 14.647 0.358 14.747 ;
    END
  END TD[1]
  PIN TD[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    ANTENNADIFFAREA 0.056 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.06 ;
    PORT
      LAYER M2 ;
        RECT 0.118 23.159 0.358 23.259 ;
    END
  END TD[2]
  PIN TD[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    ANTENNADIFFAREA 0.056 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.06 ;
    PORT
      LAYER M2 ;
        RECT 0.118 31.671 0.358 31.771 ;
    END
  END TD[3]
  PIN TD[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    ANTENNADIFFAREA 0.056 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.06 ;
    PORT
      LAYER M2 ;
        RECT 0.118 40.183 0.358 40.283 ;
    END
  END TD[4]
  PIN TD[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    ANTENNADIFFAREA 0.056 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.06 ;
    PORT
      LAYER M2 ;
        RECT 0.118 48.695 0.358 48.795 ;
    END
  END TD[5]
  PIN TD[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    ANTENNADIFFAREA 0.056 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.06 ;
    PORT
      LAYER M2 ;
        RECT 0.118 57.207 0.358 57.307 ;
    END
  END TD[6]
  PIN TD[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    ANTENNADIFFAREA 0.056 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.06 ;
    PORT
      LAYER M2 ;
        RECT 0.118 65.719 0.358 65.819 ;
    END
  END TD[7]
  PIN BWM[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    ANTENNADIFFAREA 0.056 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.06 ;
    PORT
      LAYER M2 ;
        RECT 0.118 9.396 0.358 9.496 ;
    END
  END BWM[0]
  PIN BWM[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    ANTENNADIFFAREA 0.056 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.06 ;
    PORT
      LAYER M2 ;
        RECT 0.118 17.908 0.358 18.008 ;
    END
  END BWM[1]
  PIN BWM[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    ANTENNADIFFAREA 0.056 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.06 ;
    PORT
      LAYER M2 ;
        RECT 0.118 26.42 0.358 26.52 ;
    END
  END BWM[2]
  PIN BWM[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    ANTENNADIFFAREA 0.056 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.06 ;
    PORT
      LAYER M2 ;
        RECT 0.118 34.932 0.358 35.032 ;
    END
  END BWM[3]
  PIN BWM[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    ANTENNADIFFAREA 0.056 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.06 ;
    PORT
      LAYER M2 ;
        RECT 0.118 43.444 0.358 43.544 ;
    END
  END BWM[4]
  PIN BWM[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    ANTENNADIFFAREA 0.056 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.06 ;
    PORT
      LAYER M2 ;
        RECT 0.118 51.956 0.358 52.056 ;
    END
  END BWM[5]
  PIN BWM[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    ANTENNADIFFAREA 0.056 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.06 ;
    PORT
      LAYER M2 ;
        RECT 0.118 60.468 0.358 60.568 ;
    END
  END BWM[6]
  PIN BWM[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    ANTENNADIFFAREA 0.056 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.06 ;
    PORT
      LAYER M2 ;
        RECT 0.118 68.98 0.358 69.08 ;
    END
  END BWM[7]
  PIN TBWM[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    ANTENNADIFFAREA 0.056 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.06 ;
    PORT
      LAYER M2 ;
        RECT 0.118 9.066 0.358 9.166 ;
    END
  END TBWM[0]
  PIN TBWM[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    ANTENNADIFFAREA 0.056 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.06 ;
    PORT
      LAYER M2 ;
        RECT 0.118 17.578 0.358 17.678 ;
    END
  END TBWM[1]
  PIN TBWM[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    ANTENNADIFFAREA 0.056 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.06 ;
    PORT
      LAYER M2 ;
        RECT 0.118 26.09 0.358 26.19 ;
    END
  END TBWM[2]
  PIN TBWM[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    ANTENNADIFFAREA 0.056 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.06 ;
    PORT
      LAYER M2 ;
        RECT 0.118 34.602 0.358 34.702 ;
    END
  END TBWM[3]
  PIN TBWM[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    ANTENNADIFFAREA 0.056 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.06 ;
    PORT
      LAYER M2 ;
        RECT 0.118 43.114 0.358 43.214 ;
    END
  END TBWM[4]
  PIN TBWM[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    ANTENNADIFFAREA 0.056 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.06 ;
    PORT
      LAYER M2 ;
        RECT 0.118 51.626 0.358 51.726 ;
    END
  END TBWM[5]
  PIN TBWM[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    ANTENNADIFFAREA 0.056 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.06 ;
    PORT
      LAYER M2 ;
        RECT 0.118 60.138 0.358 60.238 ;
    END
  END TBWM[6]
  PIN TBWM[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    ANTENNADIFFAREA 0.056 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.06 ;
    PORT
      LAYER M2 ;
        RECT 0.118 68.65 0.358 68.75 ;
    END
  END TBWM[7]
  PIN BADIO[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
        RECT 0.118 6.437 0.358 6.537 ;
    END
  END BADIO[0]
  PIN BADIO[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
        RECT 0.118 14.949 0.358 15.049 ;
    END
  END BADIO[1]
  PIN BADIO[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
        RECT 0.118 23.461 0.358 23.561 ;
    END
  END BADIO[2]
  PIN BADIO[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
        RECT 0.118 31.973 0.358 32.073 ;
    END
  END BADIO[3]
  PIN BADIO[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
        RECT 0.118 40.485 0.358 40.585 ;
    END
  END BADIO[4]
  PIN BADIO[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
        RECT 0.118 48.997 0.358 49.097 ;
    END
  END BADIO[5]
  PIN BADIO[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
        RECT 0.118 57.509 0.358 57.609 ;
    END
  END BADIO[6]
  PIN BADIO[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
        RECT 0.118 66.021 0.358 66.121 ;
    END
  END BADIO[7]
  PIN AWT
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    ANTENNADIFFAREA 0.056 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0536 ;
    PORT
      LAYER C1 ;
        RECT 0.118 113.186 0.358 113.286 ;
    END
  END AWT
  PIN LVTEST
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    ANTENNADIFFAREA 0.056 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0536 ;
    PORT
      LAYER C1 ;
        RECT 0.118 85.284 0.358 85.384 ;
    END
  END LVTEST
  PIN VSB400
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER C1 ;
        RECT 0.118 94.886 0.358 94.986 ;
    END
  END VSB400
  PIN VSB300
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER C1 ;
        RECT 0.118 93.976 0.358 94.076 ;
    END
  END VSB300
  PIN VSB200
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER C1 ;
        RECT 0.118 83.021 0.358 83.121 ;
    END
  END VSB200
  PIN VSB100
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER C1 ;
        RECT 0.118 78.691 0.358 78.791 ;
    END
  END VSB100
  PIN RA
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    ANTENNADIFFAREA 0.056 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0536 ;
    PORT
      LAYER M2 ;
        RECT 0.118 70.198 0.358 70.298 ;
    END
  END RA
  PIN WM[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    ANTENNADIFFAREA 0.056 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0536 ;
    PORT
      LAYER C1 ;
        RECT 0.118 99.686 0.358 99.786 ;
    END
  END WM[0]
  PIN WM[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    ANTENNADIFFAREA 0.056 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0536 ;
    PORT
      LAYER C1 ;
        RECT 0.118 101.191 0.358 101.291 ;
    END
  END WM[1]
  PIN WM[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    ANTENNADIFFAREA 0.056 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0536 ;
    PORT
      LAYER C1 ;
        RECT 0.118 102.101 0.358 102.201 ;
    END
  END WM[2]
  PIN RM[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    ANTENNADIFFAREA 0.056 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0536 ;
    PORT
      LAYER C1 ;
        RECT 0.118 104.496 0.358 104.596 ;
    END
  END RM[0]
  PIN RM[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    ANTENNADIFFAREA 0.056 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0536 ;
    PORT
      LAYER C1 ;
        RECT 0.118 105.996 0.358 106.096 ;
    END
  END RM[1]
  PIN RM[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    ANTENNADIFFAREA 0.056 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0536 ;
    PORT
      LAYER C1 ;
        RECT 0.118 108.381 0.358 108.481 ;
    END
  END RM[2]
  PIN BISTE
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    ANTENNADIFFAREA 0.056 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0536 ;
    PORT
      LAYER C1 ;
        RECT 0.118 109.286 0.358 109.386 ;
    END
  END BISTE
  PIN TCLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    ANTENNADIFFAREA 0.056 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0536 ;
    PORT
      LAYER C1 ;
        RECT 0.118 86.281 0.358 86.381 ;
    END
  END TCLK
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    SHAPE ABUTMENT ;
    ANTENNADIFFAREA 0.056 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2064 ;
    PORT
      LAYER C1 ;
        RECT 0.118 86.691 0.358 86.791 ;
    END
  END CLK
  PIN TWE
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    ANTENNADIFFAREA 0.056 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0536 ;
    PORT
      LAYER C1 ;
        RECT 0.118 73.586 0.358 73.686 ;
    END
  END TWE
  PIN WE
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    ANTENNADIFFAREA 0.056 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0536 ;
    PORT
      LAYER C1 ;
        RECT 0.118 73.314 0.358 73.414 ;
    END
  END WE
  PIN TA[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    ANTENNADIFFAREA 0.056 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0536 ;
    PORT
      LAYER C1 ;
        RECT 0.118 78.391 0.358 78.491 ;
    END
  END TA[0]
  PIN TA[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    ANTENNADIFFAREA 0.056 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0536 ;
    PORT
      LAYER C1 ;
        RECT 0.118 88.296 0.358 88.396 ;
    END
  END TA[1]
  PIN TA[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    ANTENNADIFFAREA 0.056 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0536 ;
    PORT
      LAYER C1 ;
        RECT 0.118 90.976 0.358 91.076 ;
    END
  END TA[2]
  PIN TA[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    ANTENNADIFFAREA 0.056 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0536 ;
    PORT
      LAYER C1 ;
        RECT 0.118 93.096 0.358 93.196 ;
    END
  END TA[3]
  PIN TA[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    ANTENNADIFFAREA 0.056 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0536 ;
    PORT
      LAYER C1 ;
        RECT 0.118 95.776 0.358 95.876 ;
    END
  END TA[4]
  PIN TA[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    ANTENNADIFFAREA 0.056 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0536 ;
    PORT
      LAYER C1 ;
        RECT 0.118 97.896 0.358 97.996 ;
    END
  END TA[5]
  PIN TA[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    ANTENNADIFFAREA 0.056 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0536 ;
    PORT
      LAYER C1 ;
        RECT 0.118 100.576 0.358 100.676 ;
    END
  END TA[6]
  PIN TA[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    ANTENNADIFFAREA 0.056 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0536 ;
    PORT
      LAYER C1 ;
        RECT 0.118 102.696 0.358 102.796 ;
    END
  END TA[7]
  PIN TA[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    ANTENNADIFFAREA 0.056 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0536 ;
    PORT
      LAYER C1 ;
        RECT 0.118 105.414 0.358 105.514 ;
    END
  END TA[8]
  PIN TA[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    ANTENNADIFFAREA 0.056 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0536 ;
    PORT
      LAYER C1 ;
        RECT 0.118 107.496 0.358 107.596 ;
    END
  END TA[9]
  PIN A[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    ANTENNADIFFAREA 0.056 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0536 ;
    PORT
      LAYER C1 ;
        RECT 0.118 78.096 0.358 78.196 ;
    END
  END A[0]
  PIN A[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    ANTENNADIFFAREA 0.056 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0536 ;
    PORT
      LAYER C1 ;
        RECT 0.118 88.001 0.358 88.101 ;
    END
  END A[1]
  PIN A[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    ANTENNADIFFAREA 0.056 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0536 ;
    PORT
      LAYER C1 ;
        RECT 0.118 91.291 0.358 91.391 ;
    END
  END A[2]
  PIN A[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    ANTENNADIFFAREA 0.056 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0536 ;
    PORT
      LAYER C1 ;
        RECT 0.118 92.796 0.358 92.896 ;
    END
  END A[3]
  PIN A[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    ANTENNADIFFAREA 0.056 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0536 ;
    PORT
      LAYER C1 ;
        RECT 0.118 96.091 0.358 96.191 ;
    END
  END A[4]
  PIN A[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    ANTENNADIFFAREA 0.056 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0536 ;
    PORT
      LAYER C1 ;
        RECT 0.118 97.596 0.358 97.696 ;
    END
  END A[5]
  PIN A[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    ANTENNADIFFAREA 0.056 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0536 ;
    PORT
      LAYER C1 ;
        RECT 0.118 100.891 0.358 100.991 ;
    END
  END A[6]
  PIN A[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    ANTENNADIFFAREA 0.056 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0536 ;
    PORT
      LAYER C1 ;
        RECT 0.118 102.401 0.358 102.501 ;
    END
  END A[7]
  PIN A[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    ANTENNADIFFAREA 0.056 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0536 ;
    PORT
      LAYER C1 ;
        RECT 0.118 105.696 0.358 105.796 ;
    END
  END A[8]
  PIN A[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    ANTENNADIFFAREA 0.056 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0536 ;
    PORT
      LAYER C1 ;
        RECT 0.118 107.201 0.358 107.301 ;
    END
  END A[9]
  PIN TCE
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    ANTENNADIFFAREA 0.056 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0536 ;
    PORT
      LAYER C1 ;
        RECT 0.118 83.496 0.358 83.596 ;
    END
  END TCE
  PIN CE
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    ANTENNADIFFAREA 0.056 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0536 ;
    PORT
      LAYER C1 ;
        RECT 0.118 83.256 0.358 83.356 ;
    END
  END CE
  PIN SD
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    ANTENNADIFFAREA 0.056 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0536 ;
    PORT
      LAYER C1 ;
        RECT 0.118 76.594 0.358 76.694 ;
    END
  END SD
  PIN HN
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    ANTENNADIFFAREA 0.056 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0536 ;
    PORT
      LAYER C1 ;
        RECT 0.118 75.686 0.358 75.786 ;
    END
  END HN
  PIN SL
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    ANTENNADIFFAREA 0.056 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0536 ;
    PORT
      LAYER C1 ;
        RECT 0.118 72.108 0.358 72.208 ;
    END
  END SL
  PIN SZ
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    ANTENNADIFFAREA 0.056 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0536 ;
    PORT
      LAYER C1 ;
        RECT 0.118 74.784 0.358 74.884 ;
    END
  END SZ
  PIN Q[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    ANTENNADIFFAREA 0.168 ;
    PORT
      LAYER M2 ;
        RECT 0.118 123.097 0.358 123.237 ;
    END
  END Q[8]
  PIN Q[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    ANTENNADIFFAREA 0.168 ;
    PORT
      LAYER M2 ;
        RECT 0.118 131.609 0.358 131.749 ;
    END
  END Q[9]
  PIN Q[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    ANTENNADIFFAREA 0.168 ;
    PORT
      LAYER M2 ;
        RECT 0.118 140.121 0.358 140.261 ;
    END
  END Q[10]
  PIN Q[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    ANTENNADIFFAREA 0.168 ;
    PORT
      LAYER M2 ;
        RECT 0.118 148.633 0.358 148.773 ;
    END
  END Q[11]
  PIN Q[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    ANTENNADIFFAREA 0.168 ;
    PORT
      LAYER M2 ;
        RECT 0.118 157.145 0.358 157.285 ;
    END
  END Q[12]
  PIN Q[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    ANTENNADIFFAREA 0.168 ;
    PORT
      LAYER M2 ;
        RECT 0.118 165.657 0.358 165.797 ;
    END
  END Q[13]
  PIN Q[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    ANTENNADIFFAREA 0.168 ;
    PORT
      LAYER M2 ;
        RECT 0.118 174.169 0.358 174.309 ;
    END
  END Q[14]
  PIN Q[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    ANTENNADIFFAREA 0.168 ;
    PORT
      LAYER M2 ;
        RECT 0.118 182.681 0.358 182.821 ;
    END
  END Q[15]
  PIN D[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    ANTENNADIFFAREA 0.056 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.06 ;
    PORT
      LAYER M2 ;
        RECT 0.118 121.741 0.358 121.841 ;
    END
  END D[8]
  PIN D[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    ANTENNADIFFAREA 0.056 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.06 ;
    PORT
      LAYER M2 ;
        RECT 0.118 130.253 0.358 130.353 ;
    END
  END D[9]
  PIN D[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    ANTENNADIFFAREA 0.056 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.06 ;
    PORT
      LAYER M2 ;
        RECT 0.118 138.765 0.358 138.865 ;
    END
  END D[10]
  PIN D[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    ANTENNADIFFAREA 0.056 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.06 ;
    PORT
      LAYER M2 ;
        RECT 0.118 147.277 0.358 147.377 ;
    END
  END D[11]
  PIN D[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    ANTENNADIFFAREA 0.056 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.06 ;
    PORT
      LAYER M2 ;
        RECT 0.118 155.789 0.358 155.889 ;
    END
  END D[12]
  PIN D[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    ANTENNADIFFAREA 0.056 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.06 ;
    PORT
      LAYER M2 ;
        RECT 0.118 164.301 0.358 164.401 ;
    END
  END D[13]
  PIN D[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    ANTENNADIFFAREA 0.056 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.06 ;
    PORT
      LAYER M2 ;
        RECT 0.118 172.813 0.358 172.913 ;
    END
  END D[14]
  PIN D[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    ANTENNADIFFAREA 0.056 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.06 ;
    PORT
      LAYER M2 ;
        RECT 0.118 181.325 0.358 181.425 ;
    END
  END D[15]
  PIN TD[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    ANTENNADIFFAREA 0.056 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.06 ;
    PORT
      LAYER M2 ;
        RECT 0.118 122.171 0.358 122.271 ;
    END
  END TD[8]
  PIN TD[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    ANTENNADIFFAREA 0.056 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.06 ;
    PORT
      LAYER M2 ;
        RECT 0.118 130.683 0.358 130.783 ;
    END
  END TD[9]
  PIN TD[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    ANTENNADIFFAREA 0.056 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.06 ;
    PORT
      LAYER M2 ;
        RECT 0.118 139.195 0.358 139.295 ;
    END
  END TD[10]
  PIN TD[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    ANTENNADIFFAREA 0.056 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.06 ;
    PORT
      LAYER M2 ;
        RECT 0.118 147.707 0.358 147.807 ;
    END
  END TD[11]
  PIN TD[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    ANTENNADIFFAREA 0.056 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.06 ;
    PORT
      LAYER M2 ;
        RECT 0.118 156.219 0.358 156.319 ;
    END
  END TD[12]
  PIN TD[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    ANTENNADIFFAREA 0.056 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.06 ;
    PORT
      LAYER M2 ;
        RECT 0.118 164.731 0.358 164.831 ;
    END
  END TD[13]
  PIN TD[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    ANTENNADIFFAREA 0.056 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.06 ;
    PORT
      LAYER M2 ;
        RECT 0.118 173.243 0.358 173.343 ;
    END
  END TD[14]
  PIN TD[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    ANTENNADIFFAREA 0.056 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.06 ;
    PORT
      LAYER M2 ;
        RECT 0.118 181.755 0.358 181.855 ;
    END
  END TD[15]
  PIN BWM[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    ANTENNADIFFAREA 0.056 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.06 ;
    PORT
      LAYER M2 ;
        RECT 0.118 125.432 0.358 125.532 ;
    END
  END BWM[8]
  PIN BWM[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    ANTENNADIFFAREA 0.056 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.06 ;
    PORT
      LAYER M2 ;
        RECT 0.118 133.944 0.358 134.044 ;
    END
  END BWM[9]
  PIN BWM[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    ANTENNADIFFAREA 0.056 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.06 ;
    PORT
      LAYER M2 ;
        RECT 0.118 142.456 0.358 142.556 ;
    END
  END BWM[10]
  PIN BWM[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    ANTENNADIFFAREA 0.056 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.06 ;
    PORT
      LAYER M2 ;
        RECT 0.118 150.968 0.358 151.068 ;
    END
  END BWM[11]
  PIN BWM[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    ANTENNADIFFAREA 0.056 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.06 ;
    PORT
      LAYER M2 ;
        RECT 0.118 159.48 0.358 159.58 ;
    END
  END BWM[12]
  PIN BWM[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    ANTENNADIFFAREA 0.056 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.06 ;
    PORT
      LAYER M2 ;
        RECT 0.118 167.992 0.358 168.092 ;
    END
  END BWM[13]
  PIN BWM[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    ANTENNADIFFAREA 0.056 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.06 ;
    PORT
      LAYER M2 ;
        RECT 0.118 176.504 0.358 176.604 ;
    END
  END BWM[14]
  PIN BWM[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    ANTENNADIFFAREA 0.056 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.06 ;
    PORT
      LAYER M2 ;
        RECT 0.118 185.016 0.358 185.116 ;
    END
  END BWM[15]
  PIN TBWM[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    ANTENNADIFFAREA 0.056 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.06 ;
    PORT
      LAYER M2 ;
        RECT 0.118 125.102 0.358 125.202 ;
    END
  END TBWM[8]
  PIN TBWM[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    ANTENNADIFFAREA 0.056 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.06 ;
    PORT
      LAYER M2 ;
        RECT 0.118 133.614 0.358 133.714 ;
    END
  END TBWM[9]
  PIN TBWM[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    ANTENNADIFFAREA 0.056 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.06 ;
    PORT
      LAYER M2 ;
        RECT 0.118 142.126 0.358 142.226 ;
    END
  END TBWM[10]
  PIN TBWM[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    ANTENNADIFFAREA 0.056 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.06 ;
    PORT
      LAYER M2 ;
        RECT 0.118 150.638 0.358 150.738 ;
    END
  END TBWM[11]
  PIN TBWM[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    ANTENNADIFFAREA 0.056 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.06 ;
    PORT
      LAYER M2 ;
        RECT 0.118 159.15 0.358 159.25 ;
    END
  END TBWM[12]
  PIN TBWM[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    ANTENNADIFFAREA 0.056 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.06 ;
    PORT
      LAYER M2 ;
        RECT 0.118 167.662 0.358 167.762 ;
    END
  END TBWM[13]
  PIN TBWM[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    ANTENNADIFFAREA 0.056 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.06 ;
    PORT
      LAYER M2 ;
        RECT 0.118 176.174 0.358 176.274 ;
    END
  END TBWM[14]
  PIN TBWM[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    ANTENNADIFFAREA 0.056 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.06 ;
    PORT
      LAYER M2 ;
        RECT 0.118 184.686 0.358 184.786 ;
    END
  END TBWM[15]
  PIN BADIO[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
        RECT 0.118 122.473 0.358 122.573 ;
    END
  END BADIO[8]
  PIN BADIO[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
        RECT 0.118 130.985 0.358 131.085 ;
    END
  END BADIO[9]
  PIN BADIO[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
        RECT 0.118 139.497 0.358 139.597 ;
    END
  END BADIO[10]
  PIN BADIO[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
        RECT 0.118 148.009 0.358 148.109 ;
    END
  END BADIO[11]
  PIN BADIO[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
        RECT 0.118 156.521 0.358 156.621 ;
    END
  END BADIO[12]
  PIN BADIO[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
        RECT 0.118 165.033 0.358 165.133 ;
    END
  END BADIO[13]
  PIN BADIO[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
        RECT 0.118 173.545 0.358 173.645 ;
    END
  END BADIO[14]
  PIN BADIO[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
        RECT 0.118 182.057 0.358 182.157 ;
    END
  END BADIO[15]
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER C1 ;
        RECT 0.118 190.998 89.654 191.454 ;
        RECT 0.118 186.742 89.654 187.198 ;
        RECT 0.118 182.486 89.654 182.942 ;
        RECT 0.118 178.23 89.654 178.686 ;
        RECT 0.118 173.974 89.654 174.43 ;
        RECT 0.118 169.718 89.654 170.174 ;
        RECT 0.118 165.462 89.654 165.918 ;
        RECT 0.118 161.206 89.654 161.662 ;
        RECT 0.118 156.95 89.654 157.406 ;
        RECT 0.118 152.694 89.654 153.15 ;
        RECT 0.118 148.438 89.654 148.894 ;
        RECT 0.118 144.182 89.654 144.638 ;
        RECT 0.118 139.926 89.654 140.382 ;
        RECT 0.118 135.67 89.654 136.126 ;
        RECT 0.118 131.414 89.654 131.87 ;
        RECT 0.118 127.158 89.654 127.614 ;
        RECT 0.118 122.902 89.654 123.358 ;
        RECT 0.118 118.646 89.654 119.102 ;
        RECT 0.118 99.958 89.654 100.414 ;
        RECT 0.118 109.558 89.654 110.014 ;
        RECT 0.118 95.158 89.654 95.614 ;
        RECT 0.118 80.758 89.654 81.214 ;
        RECT 0.118 78.958 89.654 79.414 ;
        RECT 0.118 74.158 89.654 74.614 ;
        RECT 0.118 75.958 89.654 76.414 ;
        RECT 0.118 71.158 89.654 71.614 ;
        RECT 0.118 93.358 89.654 93.814 ;
        RECT 0.118 98.158 89.654 98.614 ;
        RECT 0.118 88.558 89.654 89.014 ;
        RECT 0.118 90.358 89.654 90.814 ;
        RECT 0.118 102.958 89.654 103.414 ;
        RECT 0.118 107.758 89.654 108.214 ;
        RECT 0.118 104.758 89.654 105.214 ;
        RECT 0.118 112.558 89.654 113.014 ;
        RECT 0.118 114.358 89.654 114.814 ;
        RECT 0.118 85.558 89.654 86.014 ;
        RECT 0.118 83.758 89.654 84.214 ;
        RECT 0.118 66.45 89.654 66.906 ;
        RECT 0.118 62.194 89.654 62.65 ;
        RECT 0.118 57.938 89.654 58.394 ;
        RECT 0.118 53.682 89.654 54.138 ;
        RECT 0.118 49.426 89.654 49.882 ;
        RECT 0.118 45.17 89.654 45.626 ;
        RECT 0.118 40.914 89.654 41.37 ;
        RECT 0.118 36.658 89.654 37.114 ;
        RECT 0.118 32.402 89.654 32.858 ;
        RECT 0.118 28.146 89.654 28.602 ;
        RECT 0.118 23.89 89.654 24.346 ;
        RECT 0.118 19.634 89.654 20.09 ;
        RECT 0.118 15.378 89.654 15.834 ;
        RECT 0.118 11.122 89.654 11.578 ;
        RECT 0.118 6.866 89.654 7.322 ;
        RECT 0.118 2.61 89.654 3.066 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER C1 ;
        RECT 0.118 193.636 89.654 194.092 ;
        RECT 0.118 189.38 89.654 189.836 ;
        RECT 0.118 185.124 89.654 185.58 ;
        RECT 0.118 180.868 89.654 181.324 ;
        RECT 0.118 176.612 89.654 177.068 ;
        RECT 0.118 172.356 89.654 172.812 ;
        RECT 0.118 168.1 89.654 168.556 ;
        RECT 0.118 163.844 89.654 164.3 ;
        RECT 0.118 159.588 89.654 160.044 ;
        RECT 0.118 155.332 89.654 155.788 ;
        RECT 0.118 151.076 89.654 151.532 ;
        RECT 0.118 146.82 89.654 147.276 ;
        RECT 0.118 142.564 89.654 143.02 ;
        RECT 0.118 138.308 89.654 138.764 ;
        RECT 0.118 134.052 89.654 134.508 ;
        RECT 0.118 129.796 89.654 130.252 ;
        RECT 0.118 125.54 89.654 125.996 ;
        RECT 0.118 121.284 89.654 121.74 ;
        RECT 0.118 117.028 89.654 117.484 ;
      LAYER C1 ;
        RECT 0.118 101.458 89.654 101.914 ;
        RECT 0.118 111.058 89.654 111.514 ;
        RECT 0.118 96.658 89.654 97.114 ;
        RECT 0.118 82.258 89.654 82.714 ;
        RECT 0.118 77.458 89.654 77.914 ;
        RECT 0.118 72.658 89.654 73.114 ;
        RECT 0.118 91.858 89.654 92.314 ;
        RECT 0.118 87.058 89.654 87.514 ;
        RECT 0.118 106.258 89.654 106.714 ;
        RECT 0.118 115.858 89.654 116.314 ;
      LAYER C1 ;
        RECT 0.118 69.088 89.654 69.544 ;
        RECT 0.118 64.832 89.654 65.288 ;
        RECT 0.118 60.576 89.654 61.032 ;
        RECT 0.118 56.32 89.654 56.776 ;
        RECT 0.118 52.064 89.654 52.52 ;
        RECT 0.118 47.808 89.654 48.264 ;
        RECT 0.118 43.552 89.654 44.008 ;
        RECT 0.118 39.296 89.654 39.752 ;
        RECT 0.118 35.04 89.654 35.496 ;
        RECT 0.118 30.784 89.654 31.24 ;
        RECT 0.118 26.528 89.654 26.984 ;
        RECT 0.118 22.272 89.654 22.728 ;
        RECT 0.118 18.016 89.654 18.472 ;
        RECT 0.118 13.76 89.654 14.216 ;
        RECT 0.118 9.504 89.654 9.96 ;
        RECT 0.118 5.248 89.654 5.704 ;
        RECT 0.118 0.992 89.654 1.448 ;
    END
    PORT

    END
    END
    PORT
      LAYER M1 ;
        RECT 89.574 194.844 89.774 195.084 ;
      LAYER M2 ;
        RECT 0 194.984 89.774 195.084 ;
        RECT 89.574 194.844 89.774 195.084 ;
      LAYER M1 ;
        RECT 89.574 116.036 89.774 116.276 ;
      LAYER M2 ;
        RECT 0 116.036 89.774 116.136 ;
        RECT 89.574 116.036 89.774 116.276 ;
      LAYER M2 ;
        RECT 0 70.436 87.243 70.536 ;
      LAYER M1 ;
        RECT 89.574 0 89.774 0.24 ;
      LAYER M2 ;
        RECT 0 0 89.774 0.1 ;
        RECT 89.574 0 89.774 0.24 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT 0.118 0 89.654 195.084 ;
    LAYER M2 ;
      RECT 0.118 0 89.654 195.084 ;
    LAYER M3 ;
      RECT 0.118 0 89.654 195.084 ;
    LAYER C1 ;
      RECT 0.118 0 89.654 195.084 ;
    LAYER M1 ;
      RECT 0 0 0.118 1.22 ;
      RECT 0 1.22 0.118 9.732 ;
      RECT 0 9.732 0.118 18.244 ;
      RECT 0 18.244 0.118 26.756 ;
      RECT 0 26.756 0.118 35.268 ;
      RECT 0 35.268 0.118 43.78 ;
      RECT 0 43.78 0.118 52.292 ;
      RECT 0 52.292 0.118 60.804 ;
      RECT 0 60.804 0.118 69.316 ;
      RECT 0 69.316 0.118 70.536 ;
    LAYER C1 ;
      RECT 0.118 76.886 0.358 76.986 ;
      RECT 0.118 77.178 0.358 77.278 ;
      RECT 0.118 73.858 0.358 73.958 ;
      RECT 0.118 72.358 0.358 72.458 ;
      RECT 0.118 106.93 0.358 107.03 ;
      RECT 0.118 81.441 0.358 81.541 ;
      RECT 0.118 110.176 0.358 110.276 ;
      RECT 0.118 112.296 0.358 112.396 ;
      RECT 0.118 115.014 0.358 115.114 ;
      RECT 0.118 81.866 0.358 81.966 ;
      RECT 0.118 110.491 0.358 110.591 ;
      RECT 0.118 112.001 0.358 112.101 ;
      RECT 0.118 115.314 0.358 115.414 ;
    LAYER M1 ;
      RECT 0 70.486 0.118 116.126 ;
      RECT 0 116.036 0.118 117.256 ;
      RECT 0 117.256 0.118 125.768 ;
      RECT 0 125.768 0.118 134.28 ;
      RECT 0 134.28 0.118 142.792 ;
      RECT 0 142.792 0.118 151.304 ;
      RECT 0 151.304 0.118 159.816 ;
      RECT 0 159.816 0.118 168.328 ;
      RECT 0 168.328 0.118 176.84 ;
      RECT 0 176.84 0.118 185.352 ;
    LAYER M2 ;
      RECT 0.118 189.837 0.358 189.937 ;
      RECT 0.118 190.267 0.358 190.367 ;
      RECT 0.118 193.528 0.358 193.628 ;
      RECT 0.118 193.198 0.358 193.298 ;
      RECT 0.118 190.569 0.358 190.669 ;
    LAYER M1 ;
      RECT 0 185.352 0.118 193.864 ;
      RECT 0 193.864 0.118 195.084 ;
    LAYER M2 ;
      RECT 1.638 77.456 1.878 77.556 ;
      RECT 1.638 77.191 1.878 77.291 ;
      RECT 1.638 72.656 1.878 72.756 ;
      RECT 1.638 72.391 1.878 72.491 ;
    LAYER C1 ;
      RECT 1.638 106.93 1.878 107.03 ;
    LAYER M2 ;
      RECT 1.638 82.256 1.878 82.356 ;
      RECT 1.638 111.041 1.878 111.141 ;
      RECT 1.638 111.431 1.878 111.531 ;
      RECT 1.638 115.841 1.878 115.941 ;
      RECT 1.638 81.991 1.878 82.091 ;
      RECT 1.638 110.792 1.878 110.892 ;
      RECT 1.638 111.68 1.878 111.78 ;
      RECT 1.638 115.592 1.878 115.692 ;
      RECT 1.638 190.569 1.878 190.669 ;
      RECT 1.638 193.528 1.878 193.628 ;
      RECT 1.638 193.198 1.878 193.298 ;
      RECT 1.638 189.837 1.878 189.937 ;
      RECT 1.638 190.266 1.878 190.366 ;
    LAYER M1 ;
      RECT 11.523 0.05 37.852 195.034 ;
    LAYER M2 ;
      RECT 11.523 0.05 37.852 195.034 ;
    LAYER M3 ;
      RECT 11.523 0.05 37.852 195.034 ;
    LAYER C1 ;
      RECT 11.523 0.05 37.852 195.034 ;
    LAYER M1 ;
      RECT 13.495 0 13.595 0.1 ;
      RECT 17.042 0 17.142 0.1 ;
      RECT 31.579 0 31.694 0.1 ;
      RECT 13.495 70.436 13.595 70.536 ;
      RECT 17.042 70.436 17.142 70.536 ;
      RECT 31.579 70.436 31.694 70.536 ;
      RECT 13.495 116.036 13.595 116.136 ;
      RECT 17.042 116.036 17.142 116.136 ;
      RECT 31.579 116.036 31.694 116.136 ;
      RECT 13.495 194.984 13.595 195.084 ;
      RECT 17.042 194.984 17.142 195.084 ;
      RECT 31.579 194.984 31.694 195.084 ;
      RECT 37.852 0.05 89.654 195.034 ;
    LAYER M2 ;
      RECT 37.852 0.05 89.654 195.034 ;
    LAYER M3 ;
      RECT 37.852 0.05 89.654 195.034 ;
    LAYER C1 ;
      RECT 37.852 0.05 89.654 195.034 ;
    LAYER M1 ;
      RECT 89.654 0 89.774 1.296 ;
      RECT 89.654 69.214 89.774 70.536 ;
    LAYER M2 ;
      RECT 89.654 70.436 89.774 70.536 ;
    LAYER M1 ;
      RECT 89.654 69.316 89.774 116.086 ;
      RECT 89.654 116.036 89.774 117.332 ;
      RECT 89.654 193.788 89.774 195.084 ;
  END
END spram_1024x16m8b1pm2re1

END LIBRARY


