// Time-stamp: <2010-11-03 1357 ronen>
//-----------------------------------------------------------------------------
// Title         : mux2to1.v
// Project   :<project>
//-----------------------------------------------------------------------------
// File          : <filename>
// Author        : Ronen Daly
// Created       : 30-05-2010
// Last modified : 30-05-2010
//-----------------------------------------------------------------------------
// Description :
// <description>
//-----------------------------------------------------------------------------
// Copyright (c)  by <company> This model is the confidential and
// proprietary property of <company> and the possession or use of this
// file requires a written license from <company>.
//------------------------------------------------------------------------------
// Modification history :
//-----------------------------------------------------------------------------
//-------------------------------------------------------------------------------------------------
// Rev.  | Date:    | Revised By:    | Description:
//=================================================================================================
// 1.0   | <moddate>| <author>       |
//       |          |                |
//-------------------------------------------------------------------------------------------------

module mux4to1 (/*AUTOARG*/
   // Outputs
   y,
   // Inputs
   s, a3, a2, a1, a0
   );


   /*********************  DEFINE  *********************/

   /*******************  PARAMETERS  *******************/

   parameter DW = 16;


   /*********************  INPUT   *********************/
   input [1:0] s;
   input [DW-1:0] a3;
   input [DW-1:0] a2;
   input [DW-1:0] a1;
   input [DW-1:0] a0;
  
   /*********************  OUTPUT  *********************/
   output reg  [DW-1:0] y; // wired reg 
  
   /*********************  INOUT  *********************/
  
   /*********************** REGS    ********************/
  
   /*********************** COMB REGS    ********************/
   // reg stm ; // wired

   /*********************   WIRE   *********************/
  
   /*********************   AUTOSAFE    **********/
  

   /****************************************************
    **********
    **********             CODE
    **********
    ****************************************************/

   always_comb
     case (s[1:0])
       2'h0 : y[DW-1:-0] = a0[DW-1:0];
       2'h1 : y[DW-1:-0] = a1[DW-1:0];
       2'h2 : y[DW-1:-0] = a2[DW-1:0];
       2'h3 : y[DW-1:-0] = a3[DW-1:0];
       default : y[DW-1:-0] = a0[DW-1:0];
     endcase
   
   
endmodule // <modulename>



